//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.7.02Beta
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Fri May 14 19:19:08 2021

module doge_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire [27:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFEFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFEDCBACDDDEFFFFFFFFFFFFFFFFEEFFFFEFFFEDDC867BDEFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFEC93DB9AE3ADEFFFFFFFFFFFFFFFEFFFFFFFEDC92A778C5DFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFEAE9C9AB98D4BDEEEEEEDDDDDDDCDDDDEEFEDB6DAB98A7BAEFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFD68DBAAAACC9B29BCCA8543322234568BDEEC28DCAA99B84CEFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFDFCBBAAAAAAABAD37432221111112211369B58CBBBA99ADDAEFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFFFEFEA8BABABAAAABBF0022110FFFFFFF00112121FDBAAAB99AD97EFFFFFFF;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFD6A9BFBBB9ABD0010FFFFFFEEEEEEFF00010EEFCBABAAACE74DFFFFFFF;
defparam prom_inst_0.INIT_RAM_0A = 256'hFFFFFFC3B9F0EBABC0F000EEFFF0FFEEEFFFFFFFFF0EEEFCBABE0D71DFFFFFFF;
defparam prom_inst_0.INIT_RAM_0B = 256'hFFFFFFB0A9F00CADF110FEEEEEFFFFEEFFFFFFEEEFF0FEF0CCB10E60CFFFFFFF;
defparam prom_inst_0.INIT_RAM_0C = 256'hFFFFFEAE98F01C0F1010FFFFEEEEFFFFFFEEEEEEEFF0DEFEFE011071CFFFFFFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFFEAE7AFF11F10FFEFFEFEEEEEEFFFFEEEEEFFFFF0EEEEF120062CFFFFFFF;
defparam prom_inst_0.INIT_RAM_0E = 256'hFFFFFEB17AF0001FFEEFEFFFEEEEEEEEEEFFEEFFFEF01FEEEDF02F83DFFFFFFF;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFFFFC38B0F01FFEEEEFEFEEEFFEEEEEEFFFFFFFFFF1FEEEEEEFF97DFFFFFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFF98CFE10FFEEEEFFFEEE0FFFFFFEFFFFEF0FEF1FFEEEFEE1EAEFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFCBDE1FFFEFEEEF0F0F0232000FFEEFFF010102FFFEEEDF01BEFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFD1E00FFEEFFEFE02455667630FFEEF056555565300EEEE03BDFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFC3F1FEF012222258888777651FEEEEF677878A74F210FEF17DFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFEB21FEF022C640006D2A877652FFEEE067885D532206E2FE03BFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFD721F013CBAEFFEEE8C69865630FEEEF59900BFFFFD7881E029EFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFEA321F0371339FFEFFFEAA976620FEFF079F225CFFFFFF592015BEFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFE8110018994333FFFFFFE9D87510FFFE1729F3344FFFFFFED1F19DFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'hFFFFFD32001F0008334CFFFFFFF35730FFEDE0731213449FFFFF860EF3DFFFFF;
defparam prom_inst_0.INIT_RAM_19 = 256'hFFFFFB20EF1C11393339FFFFFFFAD71FFFEDEF300383442FFFFFD11EE1BEEFFF;
defparam prom_inst_0.INIT_RAM_1A = 256'hFFFFE910FF0B13444348FFFFFFF5420FFEEEE0352443348FFFFFA50DE08DEFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFD61FEE034234437FFFFFFFD001FFFEFFEF1B033337FFEFFF191EE07DEFFF;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFFDB31FEEE0011334CFFFFFFF2A20FFFFFFEEF16133ADFFFFFD2FEEE06DEFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFDA21FFEEF3D401BEFFEEE9AA31EFFF0000FE03110CEDEFE6931FEF15CEFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFEA210FFFFF22A24E664FA4B20FFFF0122220002CA8F5F929310FF014BDFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFE91100FEF001242CDDEF032FE0002345665410134521121211211113ADFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFD911000F011114566777643112356555666664333455655544334442AEFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFD8111000133333445556665555677776677776654554444443334552AEFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFD8233322333334445666666666666777778788877654444443344552AEFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFE83433333333334456777666666677787820DF015764444433345553BEFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFEA454333333343456777777777777787340111111C66444333345554BEFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFEB4444443333444567777777777777785C7622111875444333344556CEFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFC5444444334445667766667777777877C7322111B75444333334558DEFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFD7444444334456666776677777777778F1222120465444333333459DEFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFE93344443444666767766766667777678D12221186544443432342AEFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFC243443433456666767767666677766779211D866544444333344CFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFD4444444334576666877767666777667861108877554444333327DFFFFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hFFFFFE8354444434565567778876666675677871A87776765444433539EFFFFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFEB5544434345667677ED688776766778941477788FB544344445CEFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hFFFFFFD9464433345666678843E887877778955A7777834A644444539DFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFEC5444333457678777610A6988788845148788F45464344445DFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFE8254333456676777778128E322E6114C26D715585433463AEFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFFFFFFEC6443334566677777770A511100246420101D6875334557CFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFFFDB44434456666677767778645677788885377765444446CDFFFFFFFF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFFFED9354334556776777777777677777777877676533455ADFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFED83553456677777777777677777777767666553454ADEFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFFFFFFFFFED8354455667776777777777777777667776554539DFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFFFFFFFFFFFC92555566777777677777777777777667555439DFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFEC945456777766767777667766677666555349CEFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFFFFFFFFFFFFEDA43467667676677777666667777665314ADEFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFDC743567677667788777667777753236BDFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFECA645676666667777666677753469CDFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFEEEC8433345555566666543258BEFEEFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFEDB864322211122233469BDFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFEEEEDCBA8656679ACDDDEEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDCCCCDDEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFFFFFFFFFDDFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFDFFDFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFDDFDDFFFFFFFFFFFFFFFFDDFFFFFFFFFDDFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFB7FFFDDFFDFFFFFFDFFFFFFFFFFFFDFFFDFFF19FDFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFF7984A0ABFFDFFDFFFFFFFFFFFFFFFFFFFFFFFF908864FFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFF8AC6AE4A69FFFFFFFFFFFFFFFFFFFFFDFDFF360C86CE0BFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFF58C68668ECE4BDFDFB73FDDBBBBF159FFFFDB8A84846CCBFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'hFFFFFFFD0C864688668E0695DDF1555555551DBB17DDAE666666AE4FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hDFFFFFF7AE8A664666666BD555532424444533537974086648668EA9FFFFFFFF;
defparam prom_inst_1.INIT_RAM_09 = 256'hFFFFFFFF080C6682680BD37466444444444445555D84AE866668E481FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFF568036668898157266467644444444644643886886484F2ABFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFB4843F8628133646646666644444466664621A669AA811A85FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFA06453AB83175446466666664446466664645888484D331C9FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFCAC423DA75442662644444666646444666644164468151FADFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFF38E251FB48646466444444466644444446265368664A15AC1FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFD7A050F54666666464444444444444444464445A666668A8A9FFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFF7A4CA534666644444647464646244464654445A8664864B8FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFD6A85226466644527499BB35746446643339558866644873FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFDD98F5466466482579FFFDFF95464667DFDFDFFB1B948647BFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFDDF894265557557BFDDDFDFDF9644644FDFFFFF5D877764673FFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFBB322651548235262BFFFFFF9446689FFFFD6CEE0E8E9889BBFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFF3D54973AAB9FFFFD98AFFFFF9564464FFF515DFDF91C494973DFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFF9B572534EEE5FFFFFFFF8DDDF7762467FBA006DDFFFFFDA955BBFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFF7D5755C2AEEEFFFFFFFFF4DFD5544647DBAAEEEFFFFFFF4A7459FFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'hFFFDDDB555522730EE01FFFFFFF59DD5462465BA953EEE3FFFFF58768FFFFFFF;
defparam prom_inst_1.INIT_RAM_19 = 256'hFFFFD9B5245005D40EC3FFFFFFF1AF74466462DE5B2E0E7FFFFF50988BBFFFFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hFFFFD3B5463E0CEE0E21FFDFFFF3C5544444473A0E00E0FFFFFF9056875FFFFF;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFD2445540E00E0DDFFFFDF0574464464650EEE00EDFFFFFD898671FFFFF;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFB12444318EE023FFFFDFF545744644444A540ECA7FFFDFDAE6865DDFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFB324444766005FFFDFFD8457244477774475A29BFDFFF59B98665BDFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFB5544662738202BF98AA095466479775555550E4E3A2AE9976A979FFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFDB355446777333444A2D37447559FFFFFDB5775355DFF1DFD11FD99FFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'hFFFDBB5555457777BDFDDDFF755579DFFFFFFFFFF977BFDFDFFFDDDDD9BFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'hFFDD9B5B7799DFFFDFFFFFFFFDDDDFFFFFFFFFDFFFFBFFFFFFFFFFFFFBBFFFFF;
defparam prom_inst_1.INIT_RAM_22 = 256'hFFDF9B9FFFDFFFFFFFFFFFFFFFFFFFFFDFFFFFBBDFDFFFFFFFFFFFFFFB9FFFFF;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFF9FBFFFFFFFFFFFFFFFFFFFFFFFFFFDFDB37A05DFDDFFFFFFFFFFD9BFFFFF;
defparam prom_inst_1.INIT_RAM_24 = 256'hFFFFBDBFFFFFFFFFFFFFFFFFFFFFFFFFFFD7620EE0068BFFFFFFFFFFD9BFFFFF;
defparam prom_inst_1.INIT_RAM_25 = 256'hFFFFDB9FFFFFFFFFFFFFFFFFFFFFFFFFFFFD47CCCACE6BDFFFFFFFFFD7FFFFFF;
defparam prom_inst_1.INIT_RAM_26 = 256'hFFFFFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFD9492ACACE2FFFFFFFFFFFD53FFFFF;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFDFF17DFFFFFFFFFFFFFFFFFFFFFFFFFFFF24ECACEE9DFFFFFFFFFFD35FFFFF;
defparam prom_inst_1.INIT_RAM_28 = 256'hFFFFF73DFFFFFFFFFFFFDFFFFFFFFDFFFFFFD8ECAE09DFFFFFFFFFFFF9BFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hFFFFFDDFDFFDFDFFFFFFFFFFFDFDFFFFFFFDD72EC08D9FFDFFFFFFFD9FDFFFFF;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFF9FFFFFDFFDFFFFDFDFFDFFFFFFFFDFDB023BFFFDFFFFFFFFF15FFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFDFFFBFFDFFFFFFFFFDFFDBDFDDFFFFFBFFFBD4C9DDFDFFFDFFFFFFBBFFFFFF;
defparam prom_inst_1.INIT_RAM_2C = 256'hFFFFFFFF9FDFDFFFFFFFFFD4E3DFFFFFFFFFFB349FDFFD6AFFFFFFD5FFFFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFF9FFDFFFFFDFFFFFFB840BBBFDFFFBD74CDFFBB540FFFFFFDB7FFFFFFF;
defparam prom_inst_1.INIT_RAM_2E = 256'hFFFFFFDF17FFFFFFFFFFFFDB3A28BB9DDF991245FFD9C06BFFFFFF5FDDFFFFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFF9BFFFFFFFFFFDFDFB744A0C5530A202455E244BDDFFFFF9BFDFFFFFF;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFFFFFFF35DFFFFFFFFFFFFFDBFEA66666C6A4A686AC1DFFDFFF73FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFDF5FFFFFFFFFFFFFDFBD9D5B17799977B79BFDFDFFB53FFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFFFF9BBDDFFFFFFFFFFFFFFDFDBDFFFFFDBFDFDFFDFDF9D9FFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_33 = 256'hFFFFFFFFFDF59BFDFFFFFFFFFFDFFFFFFFFFFFFFFDFDFDDFFF9BBFDFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFF5BBFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFDFFDB7FFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_35 = 256'hFFFFFFFFFFFFF999FFFFFFFFFFFFFFFFFFFFFFFFFFDFFFDF9B9FFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFBB97BFFFFFDFFFFFFFFFFFFFFFFDFFDDF5DBFFDFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFBDB3DFFFFFFFFFFFDFFFFFFFFFFFFB5BFBFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFF5BD7FFDFFFFFFFFDFFFFFFFDFB3BB5FFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFB1D3BDDFFFFFFFDFFDFFFFF5BB19FFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFDFFB1B9F37BDFDDDDDDFB719BF7DFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFDFFDFFD5FD9799BB99B99BF39DFDFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFDB9753F11359DFFDFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFDDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF77FFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6EFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_04 = 256'hFFFFFFFFFFE5DC5D6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6DCCCDEFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_05 = 256'hFFFFFFFFFDC55DD5CDEFFFFFFFFFFFFFFFFFFFFF7FFFFF55555DCDFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFFFFFFFF45D55DD5DC56FFFFFFF6EEEEEE67FFFFFFF6CDD5555546FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_07 = 256'hFFFFFFFF6DDDDDDDDDD555EFEE6FFFFFFFFFF6EE7FFE45DDDD5DDDDFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_08 = 256'hFFFF7FFF45D5D5DDDDD5EE6FFFFFFFFFFFFFFFFF6EEE6DD5D5DDD54FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFE5D6EDD5DDD6EEFF7FFFFFFFFFFFFFFFFFEEEE5DD5DDD5E4FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFFFFF6D5FFE5D5DEEFFFFFFFFFFFFFFFFFFFFFFFFEEEE5DDDEE6CEFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFDD5FFE5DEEFFFFFFFFFF7FFFFFFFFFFFFFFFFEE6E5D5FFE46FFFFFFFF;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFFFFFDD5FFFDEEFFFFFFFFFFFFFFFFFFFFFFFF7FFF6EEEE6EFFFCEFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFF545FFFEEFFFF7FF7FFFFFFFFFFFFFFFFFFFFFFEEEEEFFFE4EFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFF6C5FFF6F7FF7FFFFFFFFFFFFFFFFFFFFFF7FFF6EEEEEFFE4FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFF6C6F76F777FFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEE6EECFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFF4EEEFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6EEEEEEEE5FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFF5E6FFFF77FFFFF7F7FFFF77FFFFFFFFFF7FFFE66EEEEEE6FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFFFFFEEEFFFF77F7F77FFFFFFFFF7FFFFFFFFFFFFFFF6EEEEEE6FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFFFFE6FFFFFF77777FFFFFFFFFF7FFFF77FFFFFFF765E6EEEE6FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_14 = 256'hFFFFFFFF6FFFFF7E4AADD1A45FFFFFFF7FFFFFFFF76C900982C6EE66FFFFFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hFFFFFFF7EFFFF7436FFFFF7E32FFFFFFFFFFF7FF75D7FFFF7EA36EE6FFFFFFFF;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFFFFFFEFF77F3800EFF7FFFFE3FFFF7FFFFF7FF4999EFFFFFFDB6EEEFFFFFFF;
defparam prom_inst_2.INIT_RAM_17 = 256'hFFFFFFFEFFF73BA008CFFFFFFFECFFF7FFFF77FD238804FFF7FFC4EE6FFFFFFF;
defparam prom_inst_2.INIT_RAM_18 = 256'hFFFFFFEFFFF69C428817FFFFFFFD6FF7FFFFFFF94CC8006FFFFF6AEE66FFFFFF;
defparam prom_inst_2.INIT_RAM_19 = 256'hFFFFFF6FFFF51442988EFFFFFFF7CF77FFFFF76044A010CFFFFF79EEE6FFFFFF;
defparam prom_inst_2.INIT_RAM_1A = 256'hFFFFFF6FFFFC98889816FFFFFFF6AF7FFFFFFF7A101981DFFFFFEA6EE6FFFFFF;
defparam prom_inst_2.INIT_RAM_1B = 256'hFFFFF6EFFFFF218198AFFFFFFFF1677FFFFFFF7D0081997FFFFF4B6EE6FFFFFF;
defparam prom_inst_2.INIT_RAM_1C = 256'hFFFFFEFFFFF7E100997FFFFFFF547FFFFFFFF7FF39082FFFFFFF9D6EEEEFFFFF;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFFEFFFFFF752117FFFFFFEB47F7FF7FFFF77F79947FFFFF6F66EEEEEFFFFF;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFFEFFFFFFF7FCA2C555CBA5F77FFFFFF7FFF77753B4ECB936E66EE66FFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFEFFFFFF7777FE444CD5F777F77FFFFFFFF7777FFE555EE6EFFE66EFFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hFFFFFEFFFFFF7777FFFFFFFF7777FFFFFFFFFFFFF7777FFFFFFFFFFFFF6FFFFF;
defparam prom_inst_2.INIT_RAM_21 = 256'hFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFF;
defparam prom_inst_2.INIT_RAM_22 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFF;
defparam prom_inst_2.INIT_RAM_23 = 256'hFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE54D55EFFFFFFFFFFFFFF6FFFFF;
defparam prom_inst_2.INIT_RAM_24 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE29188199CFFFFFFFFFFFFF6FFFFF;
defparam prom_inst_2.INIT_RAM_25 = 256'hFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFE4E188880BFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_2.INIT_RAM_26 = 256'hFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFF7FCE9888004FFFFFFFFFFFFF7FFFFF;
defparam prom_inst_2.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF590888806FFFFFFFFFFFF77FFFFF;
defparam prom_inst_2.INIT_RAM_28 = 256'hFFFFF77FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC88881DFFFFFFFFFFFFF6FFFFFF;
defparam prom_inst_2.INIT_RAM_29 = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB009CFFFFFFFFFFFFFFEFFFFFF;
defparam prom_inst_2.INIT_RAM_2A = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE19DFFFFFFFFFFFFFF7FFFFFFF;
defparam prom_inst_2.INIT_RAM_2B = 256'hFFFFFFFEFFFFFFFFFFF7FFFFFFFFFFFFF7FFFFE93FFFFFFFFFFFFFFFEFFFFFFF;
defparam prom_inst_2.INIT_RAM_2C = 256'hFFFFFFFEFFFFFFFFFFFF7FFD4FFFFFFFFFFFFF696FFFFF54FFFFFFFFEFFFFFFF;
defparam prom_inst_2.INIT_RAM_2D = 256'hFFFFFFFFEFFFFFFFFFF7FFFF2ADFFFFFFFFFF6A3FFFFFE24FFFFFFFEFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2E = 256'hFFFFFFFF7FFFFFFFFFFFFFFFF913EFFFFFFFE216FFFF4A2EFFFF7FFEFFFFFFFF;
defparam prom_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFEFFFFFFFFFFFFFFFF391BC66E52192C6FCB126FFFFFFF6FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_30 = 256'hFFFFFFFFF77FFFFFFFFFFFFFFFFD321111992A2999194FFFFFFFF77FFFFFFFFF;
defparam prom_inst_2.INIT_RAM_31 = 256'hFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFEEEFFFFFFFFEEFFFFFFFFF77FFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_32 = 256'hFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_33 = 256'hFFFFFFFFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_34 = 256'hFFFFFFFFFFFF76FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF67FFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_35 = 256'hFFFFFFFFFFFFFF6FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFF66FFFFFFFFFFFFFFFFFFFFFFFFFFFFE6FFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFF7E7FFFFFFFFFFFFFFFFFFFFEE7FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFF7EEEFFFFFFFFFFFFFF76E6FFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE6EE6EEE6EE66E6FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF76FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[27:0],dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 4;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_04 = 256'hFFFFFFFFFFFEDCDDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCCCCDFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_05 = 256'hFFFFFFFFFDCFFFFEBCEFFFFFFFFFFFFFFFFFFFFFFFFFFFDDFFFFDCFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_06 = 256'hFFFFFFFFFCFEFFEEFECDFFFFFFFFFEEEEEEFFFFFFFFFFBEEEFFFFCFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_07 = 256'hFFFFFFFFEEEEEEEEEEEFDDEFEEFFFFFFFFFFFFEEFFFFCFEEEEFEEECFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_08 = 256'hFFFFFFFFCFEFEFEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFEEFEFEEEFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_09 = 256'hFFFFFFFFDEFFEEFEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFEEEFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0A = 256'hFFFFFFFEDEFFFEEFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0B = 256'hFFFFFFFDDEFFFEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0C = 256'hFFFFFFFDDEFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0D = 256'hFFFFFFFEDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0E = 256'hFFFFFFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_0F = 256'hFFFFFFFECFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_10 = 256'hFFFFFFFFCFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_11 = 256'hFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFEFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFECEFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFD954AA248BFFFFFFFFFFFFFFFFFD8322226BFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_15 = 256'hFFFFFFFFEFFFFFA8EFFFFFFC75FFFFFFFFFFFFFFFA9EFFFFFC68FEFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFFFFFFEFFFFE7222CFFFFFFFD7FFFFFFFFFFFFF9112DFFFFFFC8FFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_17 = 256'hFFFFFFFEFFFF8652219FFFFFFFD8FFFFFFFFFFFB57112AFFFFFF9BFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'hFFFFFFEFFFFD2884112EFFFFFFFADFFFFFFFFFF3988122CFFFFFD6FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hFFFFFFFFFFFB2894111CFFFFFFFE9FFFFFFFFFE29942228FFFFFF3FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1A = 256'hFFFFFFFFFFFA2111112CFFFFFFFC5EFFFFFFFFF5222112BFFFFFD5FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFF5212113FFFFFFFF2DFFFFFFFFFFA221213FFFFFFA8FFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFFEFFFFFFC32211EFFFFFFFB9FFFFFFFFFFFE72215EFFFFFF4DFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFEFFFFFFFB522EFFFFFFD79FFFFFFFFFFFFFF329FFFFFFDFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFFFEFFFFFFEFE9448CCB975AFFFFFFFFFFFFFFFFA86AC9639FFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hFFFFFEFFFFFFFFFFEC9999ACEFFFFFFFFFFFFFFFFFFEECCCCCEFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_21 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_22 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDDCCDEFFFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_24 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD75666766BFFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_25 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBF9777779FFFFFFFFFFFFFEFFFFF;
defparam prom_inst_3.INIT_RAM_26 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAF777787BFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_27 = 256'hFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC5777776FFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB67776DFFFFFFFFFFFFFEFFFFFF;
defparam prom_inst_3.INIT_RAM_29 = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA776BFFFFFFFFFFFFFFEFFFFFF;
defparam prom_inst_3.INIT_RAM_2A = 256'hFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF66DFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2B = 256'hFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5AFFFFFFFFFFFFFFFEFFFFFFF;
defparam prom_inst_3.INIT_RAM_2C = 256'hFFFFFFFEFFFFFFFFFFFFFFFBBFFFFFFFFFFFFFF5EFFFFFDBFFFFFFFFEFFFFFFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hFFFFFFFFEFFFFFFFFFFFFFFF76BFFFFFFFFFFF7AFFFFFE7AFFFFFFFEFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF55AFFFFFFFFF86FFFFFD77EFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFEFFFFFFFFFFFFFFFF9568BEDDC8668BEFB868FFFFFFFFEFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDA855555688865555CFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_31 = 256'hFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_32 = 256'hFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_33 = 256'hFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_34 = 256'hFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFEEFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

endmodule //doge_rom
