/*********************************************************************************************************
 **=======================================================================================================
 ** ģ �� ��:   division
 ** ��    ��:   ʵ��ʱ�ӵķ�Ƶ, ��Ƶѡ��ϵ�����û�����
 **
 ** facter: ������ѡ��
 **   0:2400
 **   1:4800    
 **	2:9600;
 **   3:19200 
 **   4:38400
 **   5:57600    
 **	6:115200;
 **   7:230400
 **	8:384000
 **   9:460800
 **
 ** ϵ��a��Ϊǰ15�η�Ƶϵ��   
 ** ϵ��b��Ϊ��16�η�Ƶϵ����ͨ����16�ν�ǰ15�η�ƵС�����ֵ����Ƶ�ʲ��롣 
 ** a��fCLK/baudRate/16 ȡ���� b��a��16��С������(��ȥΪ������λΪ��)��
 ** �� ��:   
 **    
 **
 **=======================================================================================================
 ********************************************************************************************************/


module divider (
    clk, 
    rst, 
    factor, 
    tick_out, 
    enable
);

input               clk;                                        //  ȫ��ʱ����, (ϵͳʱ��)
input               rst;                                        //  ȫ�ָ�λ��

input               enable;                                    //  ģ��ʹ����
input   [15 : 0]    factor;                                    //  ��Ƶѡ��ϵ��
output              tick_out;                                   //  ��Ƶ���



reg     [9 : 0]    rCnt;
reg                 rPlsTick;


/********************************************************************************************************
 ** �������ʱ��ʼ���Ĵ���ֵ
 ********************************************************************************************************/
initial
begin
    rCnt <= 10'h0;
    rPlsTick <= 1'b0;
end

reg[9:0] a;
reg[9:0] b;

always@(posedge clk or posedge rst)
	if(rst) begin
		a<=10'd33;
		b<=10'd26;
	end
   else begin
		case(factor)
		0:begin       //2400
			a<=10'd651;
			b<=10'd652;
		end
		1:begin        //4800
			a<=10'd325;
			b<=10'd333;
		end
		2:begin         //9600
			a<=10'd175;  
			b<=10'd187;
		end
		3:begin        //19200
			a<=10'd81;
			b<=10'd87;
		end
		4:begin        //38400
			a<=10'd41;
			b<=10'd36;
		end
		5:begin         //57600
			a<=10'd27;
			b<=10'd29;
		end
		6:begin        //115200
			a<=10'd14;
			b<=10'd7;
		end
		7:begin        //230400
			a<=10'd7;
			b<=10'd3;
		end
		8:begin         //384000
			a<=10'd4;
			b<=10'd6;
		end
		9:begin         //460800
			a<=10'd3;
			b<=10'd9;
		end

		default:begin    //57600
			a<=10'd27;
			b<=10'd29;
		end
		endcase
	end


reg[3:0] rCountBaud;
/********************************************************************************************************
 ** ������Ƶ������, �����Ƶ�������
 ********************************************************************************************************/
always @(posedge clk or posedge rst)
begin : DIV_CNT
    if (rst) begin
        rCnt    <= 10'h0;
        rPlsTick <= 1'b0;
		  rCountBaud<=4'h0;
    end
    else 
	 if (enable) begin	 
		if(rCountBaud==4'hf)begin
			if (rCnt >= b-1'b1) begin
				rPlsTick <= 1'b1;
				rCnt    <= 10'h0;
				rCountBaud<=4'b0;
			end
			else begin
				rPlsTick <= 1'b0;
				rCnt    <= rCnt +10'h1;
			end 
		end
		else begin
			if (rCnt >= a-1) begin
				rPlsTick <= 1'b1;
				rCnt    <= 10'h0;
				rCountBaud<=rCountBaud+4'b1;
			end
			else begin
				rPlsTick <= 1'b0;
				rCnt    <= rCnt +10'h1;
			end 
	   end
    end 
    else begin 
		 rPlsTick <= 1'b0;
		 rCnt     <= 16'h0;
    end
	
end


/*
 *  ����ź�
 */
assign  tick_out = rPlsTick;

endmodule

/*********************************************************************************************************
 ** End Of File
 ********************************************************************************************************/

