//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.7.03Beta
//Part Number: GW1N-LV1QN48C6/I5
//Device: GW1N-1
//Created Time: Fri May 21 17:29:53 2021

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFEDCCBA99876654332100FEDDCBAA987665433210FFEDCCBA9887654432110F;
defparam prom_inst_0.INIT_RAM_01 = 256'h98877665443321100FEEDDCBBA998776554332110FFEDDCBBA99876654432110;
defparam prom_inst_0.INIT_RAM_02 = 256'h55444333222111000FFEEEDDCCCBBAA999887766554433221100FFEEDDCCBBAA;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFEEEEEEEEEEDDDDDDDDCCCCCCBBBBBAAAA99999888877766665;
defparam prom_inst_0.INIT_RAM_04 = 256'h6666777888899999AAAABBBBBCCCCCCDDDDDDDDEEEEEEEEEEFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hABBCCDDEEFF001122334455667788999AABBCCCDDEEEFF000111222333444555;
defparam prom_inst_0.INIT_RAM_06 = 256'h1123445667899ABBCDDEFF011233455677899ABBCDDEEF00112334456677889A;
defparam prom_inst_0.INIT_RAM_07 = 256'h0112344567889ABCCDEFF012334566789AABCDDEF00123345667899ABCCDEFF0;
defparam prom_inst_0.INIT_RAM_08 = 256'hFF0122345567889ABBCDEEF0112344567889ABBCDEFF012234566789AABCDDEF;
defparam prom_inst_0.INIT_RAM_09 = 256'h56677889AABBCDDEEF0011233455677899ABBCDDEFF01123345567889AABCDDE;
defparam prom_inst_0.INIT_RAM_0A = 256'h99AAABBBCCCDDDEEEFF00011222334455566778899AABBCCDDEEFF0011223344;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000001111111122222233333444455555666677788889;
defparam prom_inst_0.INIT_RAM_0C = 256'h8888777666655555444433333222222111111110000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h433221100FFEEDDCCBBAA99887766555443322211000FFEEEDDDCCCBBBAAA999;
defparam prom_inst_0.INIT_RAM_0E = 256'hDDCBAA98876554332110FFEDDCBBA9987765543321100FEEDDCBBAA988776654;
defparam prom_inst_0.INIT_RAM_0F = 256'hEDDCBAA987665432210FFEDCBBA9887654432110FEEDCBBA9887655432210FFE;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA998877665544332211000;
defparam prom_inst_0.INIT_RAM_21 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_22 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_23 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_24 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_25 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_26 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_27 = 256'hFEEDDCCBBAA99887766554433221100FFEEDDCCBBAA99887766554433221100F;
defparam prom_inst_0.INIT_RAM_28 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_29 = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2A = 256'h00012223445566778899AABBBCDDDEFF00112233445566678889AABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2B = 256'hF0111233345566778899AAABCCCDEEEF001122334455567778999ABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2C = 256'h00012223445566778899AABBBCDDDEFF00112233445566678889AABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2D = 256'hF0111233345566778899AAABCCCDEEEF001122334455567778999ABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2E = 256'h00012223445566778899AABBBCDDDEFF00112233444566678889AABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_2F = 256'h00111233345566778899AAABCCCDEEEF001122334455567778999ABBCCDDEEFF;
defparam prom_inst_0.INIT_RAM_30 = 256'hFFEEEEDDDDCCCCBBBBAAAA999988887777666655554444333322221111000000;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_34 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_35 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_37 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3B = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFEEEEDDDDCCCCBBBBAAAA9999888877776666555544443333222211110000FF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hAAAAAAAAAAAAAAAAAAAAAA999999999999999999998888888888888888888887;
defparam prom_inst_1.INIT_RAM_01 = 256'hDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_1.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDD;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hBBBBBBBBBBBBBBBBBBBBBBCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDD;
defparam prom_inst_1.INIT_RAM_07 = 256'h88888888888888888888899999999999999999999AAAAAAAAAAAAAAAAAAAAAAB;
defparam prom_inst_1.INIT_RAM_08 = 256'h4455555555555555555555566666666666666666666677777777777777777777;
defparam prom_inst_1.INIT_RAM_09 = 256'h2222222222222222223333333333333333333333333444444444444444444444;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000000000000000000111111111111111111111111111111111112222222222;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h2222222221111111111111111111111111111111111100000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h4444444444444444444433333333333333333333333332222222222222222222;
defparam prom_inst_1.INIT_RAM_0F = 256'h7777777777777777777666666666666666666666555555555555555555555444;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_20 = 256'h1111111111111111111111111111111000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h3333333333333333333333333333333222222222222222222222222222222221;
defparam prom_inst_1.INIT_RAM_22 = 256'h5555555555555555555555555555555444444444444444444444444444444443;
defparam prom_inst_1.INIT_RAM_23 = 256'h7777777777777777777777777777777666666666666666666666666666666665;
defparam prom_inst_1.INIT_RAM_24 = 256'h9999999999999999999999999999999888888888888888888888888888888887;
defparam prom_inst_1.INIT_RAM_25 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9;
defparam prom_inst_1.INIT_RAM_26 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCB;
defparam prom_inst_1.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEED;
defparam prom_inst_1.INIT_RAM_28 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_29 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_1.INIT_RAM_2A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_1.INIT_RAM_2B = 256'h7888888888888888888888888888888899999999999999999999999999999999;
defparam prom_inst_1.INIT_RAM_2C = 256'h6666666666666666666666666666666677777777777777777777777777777777;
defparam prom_inst_1.INIT_RAM_2D = 256'h3444444444444444444444444444444455555555555555555555555555555555;
defparam prom_inst_1.INIT_RAM_2E = 256'h2222222222222222222222222222222233333333333333333333333333333333;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000011111111111111111111111111111111;
defparam prom_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h1111111111111111111111111111111111111111111111111111111111111100;
defparam prom_inst_1.INIT_RAM_32 = 256'h2222222222222222222222222222222222222222222222222222222222222211;
defparam prom_inst_1.INIT_RAM_33 = 256'h3333333333333333333333333333333333333333333333333333333333333322;
defparam prom_inst_1.INIT_RAM_34 = 256'h4444444444444444444444444444444444444444444444444444444444444433;
defparam prom_inst_1.INIT_RAM_35 = 256'h5555555555555555555555555555555555555555555555555555555555555544;
defparam prom_inst_1.INIT_RAM_36 = 256'h6666666666666666666666666666666666666666666666666666666666666655;
defparam prom_inst_1.INIT_RAM_37 = 256'h7777777777777777777777777777777777777777777777777777777777777766;
defparam prom_inst_1.INIT_RAM_38 = 256'h8888888888888888888888888888888888888888888888888888888888888877;
defparam prom_inst_1.INIT_RAM_39 = 256'h9999999999999999999999999999999999999999999999999999999999999988;
defparam prom_inst_1.INIT_RAM_3A = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA99;
defparam prom_inst_1.INIT_RAM_3B = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBAA;
defparam prom_inst_1.INIT_RAM_3C = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBB;
defparam prom_inst_1.INIT_RAM_3D = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCC;
defparam prom_inst_1.INIT_RAM_3E = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEDD;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEE;

endmodule //Gowin_pROM
