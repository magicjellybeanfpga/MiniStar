//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.7.02Beta
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Fri May 14 20:23:46 2021

module snake_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h6D4B5CCA64CA6CCB7CED7CEF7CEF748E2A446C6D852F7D0F7CEE7D2F6CCC74EC;
defparam prom_inst_0.INIT_RAM_01 = 256'h3BA63BA643A64BA70140010000E009414B49094100E0010000E001203B264B88;
defparam prom_inst_0.INIT_RAM_02 = 256'h436653E8438712020140096109410101748E3AE7118201200981014009A14B68;
defparam prom_inst_0.INIT_RAM_03 = 256'h3AC53AE61A0201003AE72A66118309624B294B4A19C319E33AE732C7014019C3;
defparam prom_inst_0.INIT_RAM_04 = 256'h29E3092000C019E4644D2A66094221E411831183010022455BEB642C2A4500E0;
defparam prom_inst_0.INIT_RAM_05 = 256'h216208A000C0222553CB1A042245538A22252205094219E453AA53AA220500E0;
defparam prom_inst_0.INIT_RAM_06 = 256'h3183296300C02A251A2509A22244538A640D63EC222409A219C319E32A4600C0;
defparam prom_inst_0.INIT_RAM_07 = 256'h3163318300A02A46098211C309A209616C4D642D53CB32A611C21A03536A1142;
defparam prom_inst_0.INIT_RAM_08 = 256'h31633183008019A3010032C73B0711A2220419C411C311C319E30982640D1142;
defparam prom_inst_0.INIT_RAM_09 = 256'h292218E100C009212A865C0C436919C3092100E02A662AA611A2096163EC1142;
defparam prom_inst_0.INIT_RAM_0A = 256'h29A308C000C022253B0843492A6519C409422205642D4329096101214B4A1142;
defparam prom_inst_0.INIT_RAM_0B = 256'h3A6521C200E053AA1A2411C319E42A4509414B8A53AB32A6014119C3092100C0;
defparam prom_inst_0.INIT_RAM_0C = 256'h432632A5010011E219E311C34308640C012011C311A211A232865BCB118200E0;
defparam prom_inst_0.INIT_RAM_0D = 256'h32E453E93B2600E011A132C75BEC53CB00E019E319E332C76C4D5BCB00E03AE7;
defparam prom_inst_0.INIT_RAM_0E = 256'h43C73B864BE84386014000C0008000A000C000C019C211A200C000E03AE653C9;
defparam prom_inst_0.INIT_RAM_0F = 256'h338533853BA64BC73B063B063AE73AE73B074327098111C2430732A553A84367;
defparam prom_inst_0.INIT_RAM_10 = 256'h336533853B8533853B85336533653B853B85336533653B8533853B8533853365;
defparam prom_inst_0.INIT_RAM_11 = 256'h33653BA633653365338533653B85336533653B8533653385336533653BA63365;
defparam prom_inst_0.INIT_RAM_12 = 256'h3365338533853B853B853B8533653B853B8533653B853B853B85338533853365;
defparam prom_inst_0.INIT_RAM_13 = 256'h3BA633443BA600C03B85336533653B853B85336533653B8500C03BA633443BA6;
defparam prom_inst_0.INIT_RAM_14 = 256'h33653B8533653B8533653B853BA6336533653BA63B8533653B8533653B853365;
defparam prom_inst_0.INIT_RAM_15 = 256'h33653BA6336533853385338533653B853B85336533853385338533653BA63365;
defparam prom_inst_0.INIT_RAM_16 = 256'h3385336533853BA5336533853BA6336433643BA6338533653BA5338533653385;
defparam prom_inst_0.INIT_RAM_17 = 256'h3385338533853385338533852B443BA53BA52B44338533853385338533853385;
defparam prom_inst_0.INIT_RAM_18 = 256'h338533653BA5338533853385338500C03BA52B44338533853385338533853385;
defparam prom_inst_0.INIT_RAM_19 = 256'h33853BA5336533643BA533853385338533643BA6338533653BA5338533653385;
defparam prom_inst_0.INIT_RAM_1A = 256'h336533653B853B8533853B8533653B853B85336533853385338533653BA63365;
defparam prom_inst_0.INIT_RAM_1B = 256'h33653BA633653365336533653BA6336533653BA63B8533653B8533653B853365;
defparam prom_inst_0.INIT_RAM_1C = 256'h3B8533653B8500E03B85336533653B853B85336533653B8500C03BA633443BA6;
defparam prom_inst_0.INIT_RAM_1D = 256'h33853B8533653B8533653B8533653B853B8533653B853B853B85338533853365;
defparam prom_inst_0.INIT_RAM_1E = 256'h338533853B8533653BA633443B85336533653B8533653385336533653BA63365;
defparam prom_inst_0.INIT_RAM_1F = 256'h3365338533853385336533653B8533853B85336533653B8533853B8533853365;
defparam prom_inst_0.INIT_RAM_20 = 256'h3B853385338553059A05C945E105E105D125B1A7FF9DFFFFFFFFFFFFFFFE52E8;
defparam prom_inst_0.INIT_RAM_21 = 256'h43444B245B057A85B1C5D145E104E105D126FEDBFF9E00000000FFFFF7FEF7FD;
defparam prom_inst_0.INIT_RAM_22 = 256'h5AE47284A9C4C965D924E104E0E4E0E5D106FEDCFFBE00000000FFFFF7FEF7FE;
defparam prom_inst_0.INIT_RAM_23 = 256'h7A649A04D144E8E4E8E4E8E4E8E4E0E5D946B987FF3DFFBEFF9EFFBEFFFD62A7;
defparam prom_inst_0.INIT_RAM_24 = 256'hA1E4B1A4D924E8E4E8C4F0C4E8C4E8E4E0E4D104B9A7FEDCFF3DFF3C9A0699E5;
defparam prom_inst_0.INIT_RAM_25 = 256'hC165C944E104E8E4E8C4F0C4E8C4E8E4E8E4E104D926C946B9A7B986B944C9A5;
defparam prom_inst_0.INIT_RAM_26 = 256'hE104E104E8E4E8C4E8C5E8C5E8C4E8C4E8C4E8C4E0E4D8E4D925D905E104E0E4;
defparam prom_inst_0.INIT_RAM_27 = 256'hE8E4E8C4E8C4F0C4E8C5E8E5E8C5E8C4E8C4E8E4E8E4E8E4E8C4E8C4F0C4F0C4;
defparam prom_inst_0.INIT_RAM_28 = 256'hF0C4F0C4E8C4F0C4F0C5F0C5E8E4E8E4E8E4E8E3E8E4E8E4F0E4E8C4E8C4E8C4;
defparam prom_inst_0.INIT_RAM_29 = 256'hE104E0E4E8E4E8C4F0C4F0C4E8C4E8E4E8E4E104D925D125C925D166C945D125;
defparam prom_inst_0.INIT_RAM_2A = 256'hC944D144E103E8E4F0C4F0C4E8C4E8E5E8C5D105B1A7FF3DFF5EFF3EFF3D9A08;
defparam prom_inst_0.INIT_RAM_2B = 256'hA9C4B9A4D923E8E4E8C4E8C4E8C4E0E5D906B946FF3DFFBFFFBFFFDFFFBEFF9E;
defparam prom_inst_0.INIT_RAM_2C = 256'h7A649224C964E904E8E4E8E3E8E4D904B985FF1CFF7DFFDFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2D = 256'h52E57285A9C5C964D924E103E8E3D904B965FF3CFF9D00000000FFFFFFFEFFFE;
defparam prom_inst_0.INIT_RAM_2E = 256'h4345530572859205B1A5D144E0E4E8E4E125B945FF3D10000000F7FFFFFEF7FD;
defparam prom_inst_0.INIT_RAM_2F = 256'h3B8543455AE57A65A1E5C945E0E4F0C4F0C4D12699E8FF9EFFFFFFFFF7FE5308;
defparam prom_inst_0.INIT_RAM_30 = 256'h338543455305728599E5D208E1E8E9A8E9A8E1E8CA2899E5728553053B453385;
defparam prom_inst_0.INIT_RAM_31 = 256'h434553256A859AC7C268D1E7E9E8E9A8E9A8E9E8D1E7C2689AC76A8553254345;
defparam prom_inst_0.INIT_RAM_32 = 256'h52E56AA5B288D228E1E8E9E8E967F9A8F9A8E967E9E8D9E8D228B28872A552E5;
defparam prom_inst_0.INIT_RAM_33 = 256'h7A65AAC8D208E9C8E9A8E987F1A8F187F187F1A8E987E9A8E9C8D208AAA88245;
defparam prom_inst_0.INIT_RAM_34 = 256'hCA27D208E1E8E9A7E9A8F1A8E987F1A8F1A8E987E9A8E9A8E9A7E9C8D9E8D1E7;
defparam prom_inst_0.INIT_RAM_35 = 256'hF1C8E9A8E9C8E9A7F1C8E9A8E9A7F1C8F1C8E9A7E9A8F1C8E9A7F1A8F188F1A8;
defparam prom_inst_0.INIT_RAM_36 = 256'hF167F188F1A8F1A8E9A8E9A7E9C8E9A7E9A7F1C8E987E9A8E9A8F1C8E9A8E9A7;
defparam prom_inst_0.INIT_RAM_37 = 256'hF988F167F188E987E9A8E9A8F1C8E9A7F187F1A8F1A8E9A8E987E9A8E9A7E9C8;
defparam prom_inst_0.INIT_RAM_38 = 256'hE987F1C8E987E987F1C8E9A7F1A8F187F187F1A8F1A8F1A8E987F1A8E987F1C8;
defparam prom_inst_0.INIT_RAM_39 = 256'hE9C8E9A8F1C8F1C8E9A8E987E987F187F187F1C8E987F1A8F1A8F1C8F1A8E987;
defparam prom_inst_0.INIT_RAM_3A = 256'hE9A8E987E9C8E9A7E987F1C8F1A8F1A8F1A8E9A7F1A8F1C8E9A8F1A8F188F1A8;
defparam prom_inst_0.INIT_RAM_3B = 256'hDA08D9E8E9C8E9A7E9A7E9A8E987E9A7F1C8E987F1A8F1A8E9A7E9C8D9E8D1E7;
defparam prom_inst_0.INIT_RAM_3C = 256'h91E5C268E1E8F1A8E9A7E9C8E9A8E9C8E987F1C8E987E9A8E9C8D208A2C87A65;
defparam prom_inst_0.INIT_RAM_3D = 256'h6A859B08C248DA08DA08E1E8E1A7E9A7F1C8E967E9E8E1E8D228B2886AC54B05;
defparam prom_inst_0.INIT_RAM_3E = 256'h4B455B057285A2C8C268D208E1A7F1C8E9A8E9E8D1E7C2489AA76A8553253B45;
defparam prom_inst_0.INIT_RAM_3F = 256'h3B6543455305728599C5D228E1E8E9A7E9A8E1C8D20899E57285530543453385;

endmodule //snake_rom
