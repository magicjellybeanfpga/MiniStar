//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.7.02Beta
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Sat May 08 16:35:34 2021

module img_rom (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFF81FFFFFFF07FFFFFFFFFFFFFF83FFFFFFF8FFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFE03FFFFF80FFFFFFFFFFFFFFFC07FFFFFC07FFFFFFFFFFFFFF80FFFFFFE07;
defparam prom_inst_0.INIT_RAM_02 = 256'h07FFFFFFFFFFFFFFFF80FFFFE03FFFFFFFFFFFFFFFF01FFFFF01FFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFF01FFF01FFFFFFFFFFFFFFFFFE03FFF80FFFFFFFFFFFFFFFFFC07FFFC;
defparam prom_inst_0.INIT_RAM_04 = 256'hF80FFFFFFFFFFFFFFFFFFFC07FC07FFFFFFFFFFFFFFFFFF80FFE03FFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFF80E03FFFFFFFFFFFFFFFFFFFF01F01FFFFFFFFFFFFFFFFFFFE03;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000007FFE0000000000000000000007FFFFC0407FFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'h00000000003FFC0000000000000000000003FFC0000000000000000000003FFE;
defparam prom_inst_0.INIT_RAM_08 = 256'hFFC0000000000000000000003FFC0000000000000000000003FFC00000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFE03FFC001F01FFFFFFFFFFFFFE03FFC000C03FFFFFFFFFFFFFE03;
defparam prom_inst_0.INIT_RAM_0A = 256'hE03FFC00FFE03FFFFFFFFDFFFE03FFC007FC07FFFFFFFFFFFFE03FFC003F80FF;
defparam prom_inst_0.INIT_RAM_0B = 256'hC07FFFFFF0007FE03FFC03FFF80FFFFFFF800FFE03FFC01FFF01FFFFFFFC03FF;
defparam prom_inst_0.INIT_RAM_0C = 256'h03FE03FF007FFFF01FFFFFC0003FE03FF807FFFE03FFFFFE0007FE03FFC07FFF;
defparam prom_inst_0.INIT_RAM_0D = 256'hFFFFE03FFFFC0F81FE03FC007FFFFC07FFFFC0F81FE03FE007FFFF80FFFFFC07;
defparam prom_inst_0.INIT_RAM_0E = 256'hC0703FE03F0007FFFFF81FFFFC0F81FE03F0007FFFFF01FFFFC0F81FE03F8007;
defparam prom_inst_0.INIT_RAM_0F = 256'hC07FFFFC3FFFFFE0007FE03F8C07FFFFE63FFFFE0003FE03F0407FFFFFC1FFFF;
defparam prom_inst_0.INIT_RAM_10 = 256'hFFFFC03FFE03FFC07FFFF01FFFFFF801FFE03FFC07FFFF81FFFFFF0007FE03FF;
defparam prom_inst_0.INIT_RAM_11 = 256'h3FFC07FFFC003FFFFFFFFFFE03FFC07FFFC007FFFFFFFFFFE03FFC07FFFE00FF;
defparam prom_inst_0.INIT_RAM_12 = 256'h80FFFFFFFBFFE03FFC07FFF0000FFFFFFFFFFE03FFC07FFF8001FFFFFFFFFFE0;
defparam prom_inst_0.INIT_RAM_13 = 256'hFE03FFC07FF807C03FFFFFE1FFE03FFC07FFC03807FFFFFF1FFE03FFC07FFE01;
defparam prom_inst_0.INIT_RAM_14 = 256'h01FF807FFFF003FE03FFC07FF00FF00FFFFF807FE03FFC07FF00FE01FFFFFC0F;
defparam prom_inst_0.INIT_RAM_15 = 256'h000FE03FFC07F807FFC03FFFE000FE03FFC07FC03FFC03FFFF001FE03FFC07FE;
defparam prom_inst_0.INIT_RAM_16 = 256'h7E03FFFF807FF00C03E03FFC07E01FFFF00FFF80007E03FFC07F00FFFE01FFFC;
defparam prom_inst_0.INIT_RAM_17 = 256'hFC03F80603FFC07807FFFFE01FE01F00E03FFC07C03FFFFC03FE01E01E03FFC0;
defparam prom_inst_0.INIT_RAM_18 = 256'hFC0403FFFFFF80700FFC0003FFC0601FFFFFF00F807FC0203FFC0700FFFFFF00;
defparam prom_inst_0.INIT_RAM_19 = 256'hFF0007FFF8003FFC0007FFFFFFE0003FFF0003FFC0007FFFFFFC0201FFE0003F;
defparam prom_inst_0.INIT_RAM_1A = 256'h03FFC003FFFFFFFF800FFFFE003FFC001FFFFFFFF8007FFFC003FFC000FFFFFF;
defparam prom_inst_0.INIT_RAM_1B = 256'hFFFFFF07FFFFF803FFC00FFFFFFFFFE03FFFFF003FFC007FFFFFFFFC01FFFFF0;
defparam prom_inst_0.INIT_RAM_1C = 256'hFFE03FFC03FFFFFFFFFFCFFFFFFE03FFC01FFFFFFFFFF8FFFFFFC03FFC00FFFF;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFE03FFC07FFFFFFFFFFFFFFFFFE03FFC07FFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1E = 256'h00000003FFC0000000000000000000003FFC0000000000000000000003FFC07F;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000003FFC0000000000000000000003FFC00000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFE0000000000000000000007FFE0000000000000000000007FFC;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2A = 256'hFFFFFFFC00000000000007FFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFFE003FF;
defparam prom_inst_0.INIT_RAM_2B = 256'h00000000003FFFFFFFFFF000000000000003FFFFFFFFFF800000000000003FFF;
defparam prom_inst_0.INIT_RAM_2C = 256'hFFFFFFFFFFF0003FFFFFFFFFFFFFFFFFFFFC00000000000007FFFFFFFFFF8000;
defparam prom_inst_0.INIT_RAM_2D = 256'hFF07FFFFFFFFFFFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFC003FFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_30 = 256'h00000FFFFFFFFFFFFF000000000001FFFFFFFFFFFFFC00000000003FFFFFFFFF;
defparam prom_inst_0.INIT_RAM_31 = 256'hFFFFFFE0000000000007FFFFFFFFFFFE0000000000007FFFFFFFFFFFF0000000;
defparam prom_inst_0.INIT_RAM_32 = 256'hFFFFFFC07FFFFFFFFFFFC01FFFFFFFF807FFFFFFFFFFFC0000000000007FFFFF;
defparam prom_inst_0.INIT_RAM_33 = 256'hFFFFFFFFFC07FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE07FFFFFFFFFFFC07FF;
defparam prom_inst_0.INIT_RAM_34 = 256'h7FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE07FF;
defparam prom_inst_0.INIT_RAM_35 = 256'h7FFFFFFFFFFFC07FFFFF00FE07FFFFFFFFFFFC07FFFFF81FE07FFFFFFFFFFFC0;
defparam prom_inst_0.INIT_RAM_36 = 256'hFC07FFFFE007E07FFFFFFFFFFFC07FFFFE00FE07FFFFFFFFFFFC07FFFFE00FE0;
defparam prom_inst_0.INIT_RAM_37 = 256'hFE07FFFFFFFFFFFC07FFFFF00FE07FFFFFFFFFFFC07FFFFE00FE07FFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_38 = 256'hFFFFC07FF1FFFFFE07FFFFFFFFFFFC07FF9FF83FE07FFFFFFFFFFFC07FFBFF01;
defparam prom_inst_0.INIT_RAM_39 = 256'hFFFFE07FFFFFFFFFFFC07FF07FFFFE07FFFFFFFFFFFC07FF0FFFFFE07FFFFFFF;
defparam prom_inst_0.INIT_RAM_3A = 256'hFFFFFFFC07FE03FFFFE07FFFFFFFFFFFC07FE03FFFFE07FFFFFFFFFFFC07FE07;
defparam prom_inst_0.INIT_RAM_3B = 256'hC00F9FFE07FFFFFFFFFFFC07FC00FDFFE07FFFFFFFFFFFC07FC01FFFFE07FFFF;
defparam prom_inst_0.INIT_RAM_3C = 256'hFFFFFFFFFFC07F800707FE07FFFFFFFFFFFC07F80078FFE07FFFFFFFFFFFC07F;
defparam prom_inst_0.INIT_RAM_3D = 256'h07F000001FE07FFFFFFFFFFFC07F000003FE07FFFFFFFFFFFC07F800307FE07F;
defparam prom_inst_0.INIT_RAM_3E = 256'h07FFFFFFFFFFFC07E000000FE07FFFFFFFFFFFC07F000001FE07FFFFFFFFFFFC;
defparam prom_inst_0.INIT_RAM_3F = 256'hFFC07FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hFFC07FFFFFFFFFFFC07FFFFFFFFE07FFFFFFFFFFFC07FFFFFFFFE07FFFFFFFFF;
defparam prom_inst_1.INIT_RAM_01 = 256'hFFFFFC0000000000007FFFFFFFFFFFC01FFFFFFFF807FFFFFFFFFFFC07FFFFFF;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000FFFFFFFFFFFFE0000000000007FFFFFFFFFFFE0000000000007FFFFFF;
defparam prom_inst_1.INIT_RAM_03 = 256'hFFFFFFFFFC00000000007FFFFFFFFFFFFF800000000001FFFFFFFFFFFFF00000;
defparam prom_inst_1.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_06 = 256'hFFFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_07 = 256'h003FFFFFFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFE00FFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_08 = 256'hFFFF00000000000007FFFFFFFFFFF0000000000000FFFFFFFFFFFF8000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'hFE0000FFFFFFFFFFFF80000000000007FFFFFFFFFFF00000000000007FFFFFFF;
defparam prom_inst_1.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFE001FFFFFFFFFFFFFFFFFFFFFE0003FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFE00FFFFFFF;
defparam prom_inst_1.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFE00FFFFFFFFFFFFFFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFF;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFC183FFFFFFFFFFFFFFFFFFFFFC007FFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFC0FF07FFFFFFFFFFFFFFFFFFFE07C07FFFFFFFFFFFFFFFFFFFF0381FFF;
defparam prom_inst_1.INIT_RAM_11 = 256'h07FFFFFFFFFFFFFFFFFF01FF81FFFFFFFFFFFFFFFFFFFC1FF03FFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hFFFF003F81FFFF03FFFFFFFFFFFFFFFFFE0FFFF07FFFFFFFFFFFFFFFFFE07FFC;
defparam prom_inst_1.INIT_RAM_13 = 256'hFFFF040001FFFFFFF8000207FFFFE0E0003FFFFFFF8000F03FFFF80FC00FFFFF;
defparam prom_inst_1.INIT_RAM_14 = 256'hFFFFF0000003FFFFFF8000001FFFFF8000000FFFFFF0000007FFFFFE000000FF;
defparam prom_inst_1.INIT_RAM_15 = 256'h0FFFFFF80000003FFFC0000000FFFFFF80000007FFFC0000001FFFFFFC000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000060000000003FFFFE000000003FC000000007FFFFF000000007FE0000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h00001FFFF800000000000000000001FFFF800000000000000000001FFFFE0000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000FFFF000000000000000000001FFFF0000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h000000007FFE0000000000000000000007FFF000000000000000000000FFFF00;
defparam prom_inst_1.INIT_RAM_1A = 256'hC0000F80000000001F00003FFC0000000000000000000003FFE0000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h00000FFF8001FF80000F80000000003FE0001FF80000F80000000003F80001FF;
defparam prom_inst_1.INIT_RAM_1C = 256'h1FF00000F8000000003C7FC001FF00000F8000000001FFF8001FF80000F80000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000001C007F000FF00000F800000000E007E000FF00000F800000000780FE00;
defparam prom_inst_1.INIT_RAM_1E = 256'hF8007E003FFFFFE0000078001F8007F00000F8000000018001F000FF00000F80;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFE00001F8000F8007E003FFFFFE00001F8000F8007E003FFFFFE00000F8001;
defparam prom_inst_1.INIT_RAM_20 = 256'h001F0003C003FFFFFE00001F8001F8003E003FFFFFE00001F8001F8003E003FF;
defparam prom_inst_1.INIT_RAM_21 = 256'h000F80000000FE007E0003C00000F80000000FC007F0003C00000F80000001F8;
defparam prom_inst_1.INIT_RAM_22 = 256'h03FFFFC0003800000F800000003F83FC0003800000F800000007F00FE0003C00;
defparam prom_inst_1.INIT_RAM_23 = 256'h800000F8000000007FFE00003800000F800000001FFFF80003800000F8000000;
defparam prom_inst_1.INIT_RAM_24 = 256'h00000000000001800000F8000000000FF000003800000F8000000003FFC00003;
defparam prom_inst_1.INIT_RAM_25 = 256'h0018000000000000000000000001800000000000000000000000180000000000;
defparam prom_inst_1.INIT_RAM_26 = 256'h0000000000000000180000000000000000000000018000000000000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000180000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h000007FFFC000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'hF80000000000000003FFFFFFFC00000000000000000FFFFFFE00000000000000;
defparam prom_inst_1.INIT_RAM_2A = 256'h000003FFFFFFFFFC000000000000001FFFFFFFFF8000000000000000FFFFFFFF;
defparam prom_inst_1.INIT_RAM_2B = 256'hFFFFF80000018000000FFFFFFFFFFF000000100000007FFFFFFFFFF000000100;
defparam prom_inst_1.INIT_RAM_2C = 256'h38000007FFFFFFFFFFFF0000018000001FFFFFFFFFFFC0000018000001FFFFFF;
defparam prom_inst_1.INIT_RAM_2D = 256'hFFFFFFFFFC00003800001FFFFFFFFFFFFF000003800000FFFFFFFFFFFFF00000;
defparam prom_inst_1.INIT_RAM_2E = 256'h0007C0000FFFFFFFFFFFFFFE00003C00007FFFFFFFFFFFFFE00003800003FFFF;
defparam prom_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFE001FF0003FFFFFFFFFFFFFFFE000FE0000FFFFFFFFFFFFFFF0;
defparam prom_inst_1.INIT_RAM_30 = 256'hFFFE0FFFF81FFFFFFFFFFFFFFFFFC1FFFC00FFFFFFFFFFFFFFFFF007FF0007FF;
defparam prom_inst_1.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFF01FFF07FFFFFFFFFFFFFFFFFE07FFF03FFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_32 = 256'hFFFFFFFE07F03FFFFFFFFFFFFFFFFFFFC0FF81FFFFFFFFFFFFFFFFFFFC1FFC07;
defparam prom_inst_1.INIT_RAM_33 = 256'h1FFFFFFFFFFFFFFFFFFFFFC1C07FFFFFFFFFFFFFFFFFFFF03F07FFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_34 = 256'hFFFFFFFFFFFF807FFFFFFFFFFFFFFFFFFFFFE083FFFFFFFFFFFFFFFFFFFFFC08;
defparam prom_inst_1.INIT_RAM_35 = 256'h00000000000000000000000000000000000000000000000000000FFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
endmodule //img_rom
